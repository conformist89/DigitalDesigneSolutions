`include "config.vh"

module top
(
    input        clk,
    input        reset_n,
    
    input  [3:0] key_sw,
    output [3:0] led,

    output [7:0] abcdefgh,
    output [3:0] digit,

    output       buzzer,

    output       hsync,
    output       vsync,
    output [2:0] rgb
);

    assign abcdefgh  = 8'hff;
    assign digit     = 4'hf;
    assign buzzer    = 1'b0;
    assign hsync     = 1'b1;
    assign vsync     = 1'b1;
    assign rgb       = 3'b0;

    wire a = ~ key_sw [0];
    wire b = ~ key_sw [1];
    
    wire result = a ^ b;

    assign led [0] = ~ result;
    
    assign led [1] = ~ (~ key_sw [0] ^ ~ key_sw [1]);

    // Exercise 1: Change the code below.
    // Assign to led [2] the result of AND operation
    
	 wire c = key_sw[2];
	 wire d = key_sw[3];
	 
	 wire result1 = c & d;
	 wire result2 = ( ~c&d ^ (d&(~c)));
//	 
	 assign led[2] =  result1;
	 assign led[3] = result2;
	 
//    assign led [2] = 1'b0;
//
//    // Exercise 2: Change the code below.
//    // Assign to led [3] the result of XOR operation
//    // without using "^" operation.
//    // Use only operations "&", "|", "~" and parenthesis, "(" and ")".
//
//    assign led [3] = 1'b0;
//	assign led = key_sw + 4'b0001;

endmodule
